/*
Van der Corput Sequence Generator (32-bit)

This SystemVerilog module implements a Van der Corput sequence generator for bases 2, 3, and 7.
The Van der Corput sequence is a low-discrepancy sequence that provides well-distributed
points in the interval [0, 1]. This implementation generates 32-bit integer outputs
scaled by base^scale.

The algorithm works by:
1. Converting the input integer k to the specified base representation
2. Reversing the digits of the base representation
3. Scaling the result by base^scale

This implementation supports:
- Base 2: Binary Van der Corput sequence
- Base 3: Ternary Van der Corput sequence  
- Base 7: Septenary Van der Corput sequence
- 32-bit integer arithmetic
- Configurable scale parameter (default 16)
*/

module vdcorput_32bit #(
    parameter BASE = 2,      // Base of the sequence (2, 3, or 7)
    parameter SCALE = 16     // Scale factor (number of digits)
) (
    input  wire        clk,           // Clock signal
    input  wire        rst_n,         // Active-low reset
    input  wire        pop_enable,    // Enable pop operation
    input  wire [31:0] seed,          // Seed value for reseed
    input  wire        reseed_enable, // Enable reseed operation
    output reg  [31:0] vdc_out,       // Van der Corput output
    output reg         valid          // Output valid flag
);

    // Internal registers
    reg [31:0] count;
    reg [31:0] factor;
    
    // Pre-computed factor values for common base/scale combinations
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            if (BASE == 2 && SCALE == 16) begin
                factor <= 32'd65536;
            end else if (BASE == 2 && SCALE == 10) begin
                factor <= 32'd1024;
            end else if (BASE == 2 && SCALE == 11) begin
                factor <= 32'd2048;
            end else if (BASE == 3 && SCALE == 16) begin
                factor <= 32'd43046721;
            end else if (BASE == 3 && SCALE == 7) begin
                factor <= 32'd2187;
            end else if (BASE == 7 && SCALE == 16) begin
                factor <= 32'd3323293056;  // Truncated to 32 bits
            end else begin
                factor <= 32'd65536;  // Default to 2^16
            end
        end
    end
    
    // Main sequential logic
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            count <= 32'd0;
            vdc_out <= 32'd0;
            valid <= 1'b0;
        end else begin
            // Handle reseed operation
            if (reseed_enable) begin
                count <= seed;
                vdc_out <= 32'd0;
                valid <= 1'b0;
            end 
            // Handle pop operation
            else if (pop_enable) begin
                count <= count + 1'b1;
                vdc_out <= calculate_vdc(count + 1'b1);
                valid <= 1'b1;
            end else begin
                valid <= 1'b0;
            end
        end
    end
    
    // Van der Corput calculation
    function [31:0] calculate_vdc;
        input [31:0] k;
        reg [31:0] k_temp;
        reg [31:0] vdc_val;
        reg [31:0] factor_temp;
        reg [31:0] remainder;
        begin
            k_temp = k;
            vdc_val = 32'd0;
            factor_temp = factor;
            
            while (k_temp != 0) begin
                factor_temp = factor_temp / BASE;
                remainder = k_temp % BASE;
                k_temp = k_temp / BASE;
                vdc_val = vdc_val + (remainder * factor_temp);
            end
            
            calculate_vdc = vdc_val;
        end
    endfunction

endmodule